----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:53:12 05/17/2022 
-- Design Name: 
-- Module Name:    ShiftModule - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ShiftModule is
port(
		a: in std_logic_vector(31 downto 0);
		y: out std_logic_vector(31 downto 0)
		);
end ShiftModule;

architecture Behavioral of ShiftModule is

	begin
	
	y <= std_logic_vector(shift_left(unsigned(a), 2));


end Behavioral;

