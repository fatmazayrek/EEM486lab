--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   21:30:19 05/08/2022
-- Design Name:   
-- Module Name:   C:/Users/Fatma/Desktop/KODLAR/Xilinx/LAB_4/Regfile_test.vhd
-- Project Name:  LAB_4
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Regfile
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY Regfile_test IS
END Regfile_test;
 
ARCHITECTURE behavior OF Regfile_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Regfile
    PORT(
         clk : IN  std_logic;
         aa : IN  std_logic_vector(4 downto 0);
         ab : IN  std_logic_vector(4 downto 0);
         aw : IN  std_logic_vector(4 downto 0);
         wren : IN  std_logic;
         wdata : IN  std_logic_vector(31 downto 0);
         a : OUT  std_logic_vector(31 downto 0);
         b : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal aa : std_logic_vector(4 downto 0) := (others => '0');
   signal ab : std_logic_vector(4 downto 0) := (others => '0');
   signal aw : std_logic_vector(4 downto 0) := (others => '0');
   signal wren : std_logic := '0';
   signal wdata : std_logic_vector(31 downto 0) := (others => '0');

 	--Outputs
   signal a : std_logic_vector(31 downto 0);
   signal b : std_logic_vector(31 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Regfile PORT MAP (
          clk => clk,
          aa => aa,
          ab => ab,
          aw => aw,
          wren => wren,
          wdata => wdata,
          a => a,
          b => b
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 10 ns;
		
		aa <= "00001";
		ab <= "01100";
		aw <= "01000";
		wren <= '0';
		wdata <= "00110010110100010010010011010010";

      wait for clk_period*5;

		aa <= "00100";
		ab <= "01100";
		aw <= "01000";
		wren <= '1';
		wdata <= "00110010110100010010010011010010";		
		
		wait for clk_period*3;

		aa <= "01000";
		ab <= "00001";
		aw <= "01000";
		wren <= '0';
		wdata <= "00110010110100010010010011010010";	
		
		wait for clk_period*3;

		--aa <= "00100";
		--ab <= "01100";
		aw <= "01100";
		wren <= '1';
		wdata <= "00110010110101010011010011011010";	
		
		wait for clk_period*3;  

		aa <= "01100";
		ab <= "00001";
		aw <= "01000";
		wren <= '0';
		wdata <= "00110010110101010011010011011010";	

      -- insert stimulus here 

      wait;
   end process;

END;
